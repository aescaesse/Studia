* C:\Users\laboratorium\Desktop\lab 2\Lab_2_1.sch

* Schematics Version 9.1 - Web Update 1
* Fri Mar 08 08:17:44 2019



** Analysis setup **
.ac DEC 10 0.001 1MEG
.OPTIONS NOBIAS
.OPTIONS NOPAGE
.OP 


* From [PSPICE NETLIST] section of pspiceev.ini:
.lib "nom.lib"

.INC "Lab_2_1.net"
.INC "Lab_2_1.als"


.probe


.END
