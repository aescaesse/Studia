* C:\Users\laboratorium\Desktop\lab 2\lab 2.3\lab 2.3.sch

* Schematics Version 9.1 - Web Update 1
* Fri Mar 08 08:49:08 2019



** Analysis setup **
.ac DEC 10 0.001 1MEG
.OPTIONS NOBIAS
.OPTIONS NOPAGE
.OP 


* From [PSPICE NETLIST] section of pspiceev.ini:
.lib "nom.lib"

.INC "lab 2.3.net"
.INC "lab 2.3.als"


.probe


.END
