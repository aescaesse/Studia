* C:\Users\laboratorium\Desktop\lab2.3.sch

* Schematics Version 9.1 - Web Update 1
* Fri Mar 01 08:55:36 2019



** Analysis setup **
.tran 10m 500m
.OPTIONS NOBIAS
.OPTIONS NOPAGE
.OP 


* From [PSPICE NETLIST] section of pspiceev.ini:
.lib "nom.lib"

.INC "lab2.3.net"
.INC "lab2.3.als"


.probe


.END
